


package RISCV_pkg;


 import uvm_pkg::*;
 
 `include "uvm_macros.svh"
  

  `include "RISCV_seq_item.sv"
  `include "Sequence.sv"
  `include "Sequencer.sv"   
  `include "Driver.sv"  
  `include "Monitor.sv"
  `include "Coverage_collector.sv"
  `include "Agent.sv"  
  `include "Environment.sv"  
  `include "RISCV_Test.sv"

 

endpackage 

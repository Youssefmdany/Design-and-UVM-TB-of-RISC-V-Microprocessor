


package RISCV_pkg;


 import uvm_pkg::*;
 
 `include "uvm_macros.svh"
  
  `include "mem_ref_model.sv" 
  `include "reg_ref_model.sv" 
  `include "RISCV_seq_item.sv"
  `include "Sequence.sv"
  `include "Sequencer.sv"   
  `include "Driver.sv"  
  `include "Monitor.sv"
  `include "Coverage_collector.sv"
  `include "Agent.sv" 
  `include "Scoreboard.sv"   
  `include "Environment.sv"  
  `include "RISCV_Test.sv"



endpackage 
